//basic decryption and

module basic_and (
	input logic a_i, b_i, 
	output c_o
	);
  assign c_o = a_i & b_i;
  endmodule
