//basic decryption and
module basic_and (input wire in_a, in_b, output out_c);
  assign out_c = in_a & in_b;
